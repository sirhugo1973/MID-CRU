-- ram_s3.vhd

-- Generated using ACDS version 19.1 240

library IEEE;
library ram_1port_191;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ram_s3 is
	port (
		data    : in  std_logic_vector(63 downto 0) := (others => '0'); --    data.datain
		q       : out std_logic_vector(63 downto 0);                    --       q.dataout
		address : in  std_logic_vector(7 downto 0)  := (others => '0'); -- address.address
		wren    : in  std_logic                     := '0';             --    wren.wren
		clock   : in  std_logic                     := '0';             --   clock.clk
		rden    : in  std_logic                     := '0'              --    rden.rden
	);
end entity ram_s3;

architecture rtl of ram_s3 is
	component ram_s3_ram_1port_191_ef7qrwa_cmp is
		port (
			data    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- datain
			q       : out std_logic_vector(63 downto 0);                    -- dataout
			address : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			wren    : in  std_logic                     := 'X';             -- wren
			clock   : in  std_logic                     := 'X';             -- clk
			rden    : in  std_logic                     := 'X'              -- rden
		);
	end component ram_s3_ram_1port_191_ef7qrwa_cmp;

	for ram_1port_0 : ram_s3_ram_1port_191_ef7qrwa_cmp
		use entity ram_1port_191.ram_s3_ram_1port_191_ef7qrwa;
begin

	ram_1port_0 : component ram_s3_ram_1port_191_ef7qrwa_cmp
		port map (
			data    => data,    --    data.datain
			q       => q,       --       q.dataout
			address => address, -- address.address
			wren    => wren,    --    wren.wren
			clock   => clock,   --   clock.clk
			rden    => rden     --    rden.rden
		);

end architecture rtl; -- of ram_s3
