-------------------------------------------------------------------------------
-- --
-- University of Cape Town, Electrical Engineering Department--
-- --
-------------------------------------------------------------------------------
--
-- unit name: o2_h_synth.vhd
--
-- author: Nathan Boyles (nathanh.boyles@gmail.com)
--
-- date: 07/04/2020
--
-- version: 0.1
--
-- description: Synthesizes O2 header from local and regional card ID
--
-- dependencies: var_defs_pkg.vhd; util_pkg.vhd; sig_defs_pkg.vhd;
--
-- references: <reference one>
-- <reference two> ...
--
-- modified by: Nathan Boyles (nathanh.boyles@gmail.com)
--
-------------------------------------------------------------------------------
-- last changes: 07/04/2020 NB Full System Integration
-- <extended description>
-------------------------------------------------------------------------------
-- TODO: <next thing to do>
-- <another thing to do>
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.sig_defs_pkg.all;
use work.util_pkg.all;
use work.var_defs_pkg.all;

--=============================================================================
--Entity declaration for o2_h_synth
--=============================================================================
entity o2_h_synth is
port(
	--global input signals
	clk_i: in std_logic; --local bus clock
	reset_n_i: in std_logic; --reset =0: reset active
									 --      =1: no reset
	o2_h_synthI: in t_o2_h_synthI; --GBT data signals defined in sig_defs_pkg
	
	--global output signals
	o2_h_synthO: out t_o2_h_synthO
);
end entity o2_h_synth;

--===============================================================================
--Architecture declaration
--===============================================================================

architecture behaviour of o2_h_synth is

	--===============================================================================
	--Signal Aliasing
	--===============================================================================
	
	--===============================================================================
	--Signal Declaration
	--===============================================================================
	
	--===============================================================================
	--Component Declaration
	--===============================================================================
	
	--===============================================================================
	--Component Instantiation
	--===============================================================================
	
	--===============================================================================
	--Architecture begin
	--===============================================================================
begin

process(clk_i,o2_h_synthI.o2_h_synth_valid_i) is
	variable id: std_logic_vector(7 downto 0);
	begin
		if rising_edge(clk_i) then
			if o2_h_synthI.o2_h_synth_valid_i='1' then
				id:=o2_h_synthI.o2_h_synth_reg_id_i & o2_h_synthI.o2_h_synth_loc_id_i;
				
				case id is 
					when x"00" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100100000000001";
					when x"01" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101100000000001";
					when x"02" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101100000000010";
					when x"03" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110100000000001";
					when x"04" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110100000000010";
					when x"05" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111100000000001";
					when x"06" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111100000000010";
					when x"07" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001100000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011100000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101100000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111100000000100";
					when x"08" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111100000000001";
					when x"09" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111100000000010";
					when x"0A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001100000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011100000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101100000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111100000000100";
					when x"0B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000100000000001";
					when x"0C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000100000000010";
					when x"0D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001100000000001";
					when x"0E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001100000000010";
					when x"0F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010100000000001";
					when x"10" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000000010";
					when x"11" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000000100";
					when x"12" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000001000";
					when x"13" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000010000000001";
					when x"14" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000010000000010";
					when x"15" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001010000000001";
					when x"16" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001010000000010";
					when x"17" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010010000000001";
					when x"18" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000000010";
					when x"19" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000000100";
					when x"1A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001010000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011010000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101010000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111010000001000";
					when x"1B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000010000000001";
					when x"1C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000010000000010";
					when x"1D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001010000000001";
					when x"1E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001010000000010";
					when x"1F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010010000000001";
					when x"20" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100001000000001";
					when x"21" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101001000000001";
					when x"22" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101001000000010";
					when x"23" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110001000000001";
					when x"24" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110001000000010";
					when x"25" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111001000000001";
					when x"26" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111001000000010";
					when x"27" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001001000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011001000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101001000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111001000000100";
					when x"28" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001001000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011001000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101001000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111001000001000";
					when x"29" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110001000000001";
					when x"2A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110001000000010";
					when x"2B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000001000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010001000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100001000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110001000000100";
					when x"2C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000001000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010001000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100001000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110001000001000";
					when x"2D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111001000000001";
					when x"30" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100000100000001";
					when x"31" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000100000001";
					when x"32" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000100000010";
					when x"33" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000100000001";
					when x"34" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000100000010";
					when x"35" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000100000001";
					when x"36" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000100000010";
					when x"37" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000100000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000100000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000100000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000100000100";
					when x"38" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000100001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000100001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000100001000";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000100001000";
					when x"39" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000100000001";
					when x"3A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000100000010";
					when x"3B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000100000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000100000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000100000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000100000100";
					when x"3C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000100001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000100001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000100001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000100001000";
					when x"3D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000100000001";
					when x"40" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100000010000001";
					when x"41" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000010000001";
					when x"42" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000010000010";
					when x"43" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000010000001"; 
					when x"44" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000010000010";
					when x"45" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000010000001";
					when x"46" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000010000010";
					when x"47" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000010000001";
					when x"48" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000010000010";
					when x"49" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000010000001";
					when x"4A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000010000010";
					when x"4B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000010000001";
					when x"4C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000010000010";
					when x"4D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000010000001";
					when x"4E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000010000010";
					when x"4F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010000010000001";
					when x"50" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100000001000001";
					when x"51" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000001000001";
					when x"52" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000001000010";
					when x"53" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000001000001";
					when x"54" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000001000010";
					when x"55" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000001000001";
					when x"56" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000001000010";
					when x"57" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000001000001";
					when x"58" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000001000010";
					when x"59" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000001000001";
					when x"5A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000001000010";
					when x"5B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000001000001";
					when x"5C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000001000010";
					when x"5D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000001000001";
					when x"5E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000001000010";
					when x"5F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010000001000001";
					when x"60" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100000000100001";
					when x"61" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000000100001";
					when x"62" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000000100010";
					when x"63" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000000100001";
					when x"64" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000000100010";
					when x"65" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000000100001";
					when x"66" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000000100010";
					when x"67" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000000100001";
					when x"68" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000000100010";
					when x"69" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000000100001";
					when x"6A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000000100010";
					when x"6B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000000100001";
					when x"6C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000000100010";
					when x"6D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000000100001";
					when x"6E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000000100010";
					when x"6F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010000000100001";
					when x"70" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001110000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100000000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110010000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000100000000010001";
					when x"71" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001111000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100001000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110011000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000101000000010001";
					when x"72" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010000000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100010000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110100000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000110000000010001";
					when x"73" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0010001000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0100011000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110101000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000111000000010001";
					when x"74" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010010000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100100000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110110000000010001";
					when x"75" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000001000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010011000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100101000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0110111000000010001";
					when x"76" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000010000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010100000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100110000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111000000000010001";
					when x"77" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000011000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010101000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0100111000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111001000000010001";
					when x"78" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000100000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010110000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101000000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111010000000010001";
					when x"80" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011100000000001";
					when x"81" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010100000000001";
					when x"82" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010100000000010";
					when x"83" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001100000000001";
					when x"84" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001100000000010";
					when x"85" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000100000000001";
					when x"86" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000100000000010";
					when x"87" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010100000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100100000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110100000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000100000000100";
					when x"88" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110100000000001";
					when x"89" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110100000000010";
					when x"8A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000100000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010100000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100100000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110100000000100";
					when x"8B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101100000000001";
					when x"8C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101100000000010";
					when x"8D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100100000000001";
					when x"8E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110100000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000100000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010100000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100100000000010";
					when x"8F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101100000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111100000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001100000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011100000000001";
					when x"90" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000000010";
					when x"91" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000000100";
					when x"92" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000001000";
					when x"93" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101010000000001";
					when x"94" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101010000000010";
					when x"95" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100010000000001";
					when x"96" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100010000000010";
					when x"97" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011010000000001";
					when x"98" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000000010";
					when x"99" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000000100";
					when x"9A" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000010000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010010000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100010000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110010000001000";
					when x"9B" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101010000000001";
					when x"9C" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101010000000010";
					when x"9D" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100010000000001";
					when x"9E" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110010000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000010000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010010000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100010000000010";
					when x"9F" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101010000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111010000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001010000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011010000000001";
					when x"A0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011001000000001";
					when x"A1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010001000000001";
					when x"A2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010001000000010";
					when x"A3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001001000000001";
					when x"A4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001001000000010";
					when x"A5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000001000000001";
					when x"A6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000001000000010";
					when x"A7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010001000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100001000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110001000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000001000000100";
					when x"A8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010001000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100001000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110001000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000001000001000";
					when x"A9" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111001000000001";
					when x"AA" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001001000000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011001000000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101001000000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111001000000010";
					when x"AB" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001001000000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011001000000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101001000000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111001000000100";
					when x"AC" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001001000001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011001000001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101001000001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111001000001000";
					when x"AD" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000001000000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010001000000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100001000000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110001000000001";
					when x"B0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011000100000001";
					when x"B1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000100000001";
					when x"B2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000100000010";
					when x"B3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000100000001";
					when x"B4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000100000010";
					when x"B5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000100000001";
					when x"B6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000100000010";
					when x"B7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000100000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000100000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000100000100";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000100000100";
					when x"B8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000100001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000100001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000100001000";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000100001000";
					when x"B9" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000100000001";
					when x"BA" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000100000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000100000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000100000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000100000010";
					when x"BB" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000100000100";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000100000100";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000100000100";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000100000100";
					when x"BC" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000100001000";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000100001000";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000100001000";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000100001000";
					when x"BD" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000100000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000100000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000100000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000100000001";
					when x"C0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011000010000001";
					when x"C1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000010000001";
					when x"C2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000010000010";
					when x"C3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000010000001";
					when x"C4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000010000010";
					when x"C5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000010000001";
					when x"C6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000010000010";
					when x"C7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000010000001";
					when x"C8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000010000010";
					when x"C9" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000010000001";
					when x"CA" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000010000010";
					when x"CB" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000010000001";
					when x"CC" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000010000010";
					when x"CD" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000010000001";
					when x"CE" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000010000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000010000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000010000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000010000010";
					when x"CF" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101000010000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111000010000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001000010000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011000010000001";
					when x"D0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011000001000001";
					when x"D1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000001000001";
					when x"D2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000001000010";
					when x"D3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000001000001";
					when x"D4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000001000010";
					when x"D5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000001000001";
					when x"D6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000001000010";
					when x"D7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000001000001";
					when x"D8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000001000010";
					when x"D9" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000001000001";
					when x"DA" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000001000010";
					when x"DB" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000001000001";
					when x"DC" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000001000010";
					when x"DD" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000001000001";
					when x"DE" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000001000010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000001000010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000001000010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000001000010";
					when x"DF" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101000001000001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111000001000001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001000001000001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011000001000001";
					when x"E0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011000000100001";
					when x"E1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000000100001";
					when x"E2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000000100010";
					when x"E3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000000100001";
					when x"E4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000000100010";
					when x"E5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000000100001";
					when x"E6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000000100010";
					when x"E7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000000100001";
					when x"E8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000000100010";
					when x"E9" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000000100001";
					when x"EA" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000000100010";
					when x"EB" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000000100001";
					when x"EC" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000000100010";
					when x"ED" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000000100001";
					when x"EE" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000000100010";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000000100010";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000000100010";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000000100010";
					when x"EF" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101000000100001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111000000100001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001000000100001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011000000100001";
					when x"F0" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001101000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011111000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110001000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000011000000010001";
					when x"F1" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001100000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011110000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0110000000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000010000000010001";
					when x"F2" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001011000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011101000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101111000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000001000000010001";
					when x"F3" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001010000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011100000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101110000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="1000000000000010001";
					when x"F4" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001001000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011011000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101101000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111111000000010001";
					when x"F5" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0001000000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011010000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101100000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111110000000010001";
					when x"F6" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000111000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011001000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101011000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111101000000010001";
					when x"F7" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000110000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0011000000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101010000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111100000000010001";
					when x"F8" =>
							o2_h_synthO.o2_h_synth_mt11_o<="0000101000000010001";
							o2_h_synthO.o2_h_synth_mt12_o<="0010111000000010001";
							o2_h_synthO.o2_h_synth_mt21_o<="0101001000000010001";
							o2_h_synthO.o2_h_synth_mt22_o<="0111011000000010001";
					when others=>
							o2_h_synthO.o2_h_synth_mt11_o<="0000000000000000000";
							o2_h_synthO.o2_h_synth_mt12_o<="0000000000000000000";
							o2_h_synthO.o2_h_synth_mt21_o<="0000000000000000000";
							o2_h_synthO.o2_h_synth_mt22_o<="0000000000000000000";
				end case;
				o2_h_synthO.o2_h_synth_valid_o<='1';
			elsif o2_h_synthI.o2_h_synth_valid_i='0' then
				o2_h_synthO.o2_h_synth_valid_o<='0';
			end if;
		end if;
	end process;

end architecture behaviour;
--===============================================================================
--Architecture end
--===============================================================================