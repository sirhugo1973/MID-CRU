-------------------------------------------------------------------------------
-- --
-- University of Cape Town, Electrical Engineering Department--
-- --
-------------------------------------------------------------------------------
--
-- unit name: s2_pipe.vhd
--
-- author: Nathan Boyles (nathanh.boyles@gmail.com
--
-- date: $Date: 07/04/2020
--
-- version: 0.1
--
-- description: Stage 3 Pipeline module
--
-- dependencies: <entity name>, ...
--
-- references: <reference one>
-- <reference two> ...
--
-- modified by: Nathan Boyles (nathanh.boyles@gmail.com)
--
-------------------------------------------------------------------------------
-- last changes: 07/04/2020 NB Full System Integration
-- <extended description>
-------------------------------------------------------------------------------
-- TODO: <next thing to do>
-- <another thing to do>
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.sig_defs_pkg.all;
use work.util_pkg.all;
use work.var_defs_pkg.all;

entity s3_pipe is
port(clk_i: in std_logic;
	  reset_n_i: in std_logic;
	  s3_pipeI: in t_s2_pipeO;
	  s3_busy_o: out std_logic;
	  s3_pipeO: out t_s3_pipeO
);
end entity s3_pipe;

architecture main of s3_pipe is

	--===========================================================================
	--Signal Declaration
	--===========================================================================
	
	type data_port_arr_i is array (0 to 3) of std_logic_vector(63 downto 0);
	signal s_data_port_arr_i: data_port_arr_i := (others => x"0000000000000000");
	
	type data_port_arr_o is array (0 to 3) of std_logic_vector(63 downto 0);
	signal s_data_port_arr_o: data_port_arr_o;--:= (others => x"0000000000000000");
	
	type addr_port_arr_i is array (0 to 3) of std_logic_vector(7 downto 0);
	signal s_addr_port_arr_i: addr_port_arr_i:=(others =>"00000000");
	
	
	signal s3_pipe_rden_i: std_logic_vector(3 downto 0):=x"0";
	signal s3_pipe_wren_i: std_logic_vector(3 downto 0):=x"0";

	--===========================================================================
	--Component Declaration
	--===========================================================================
	 component ram_s3 is
        port (
            data    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- datain
            q       : out std_logic_vector(63 downto 0);                    -- dataout
            address : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
            wren    : in  std_logic                     := 'X';             -- wren
            clock   : in  std_logic                     := 'X';             -- clk
            rden    : in  std_logic                     := 'X'              -- rden
        );
	 end component ram_s3;

	 --==========================================================================
	 --Component Instatiation
	 --==========================================================================
	 begin
	 
	 s_ram: for i in 3 downto 0 generate
	
	 begin
	 u0 : component ram_s3
				port map (
            data    => s_data_port_arr_i(i),    --    data.datain
            q       => s_data_port_arr_o(i),       --       q.dataout
            address => s_addr_port_arr_i(i), -- address.address
            wren    => s3_pipe_wren_i(i),    --    wren.wren
            clock   => clk_i,    --   clock.clk
				rden    => s3_pipe_rden_i(i)     --    rden.rden
			);
	end generate s_ram;
	
	process(clk_i,reset_n_i,s3_pipeI) is
	
		variable s3_flag: integer range 0 to 129:=0;
		variable s3_pipe_v: t_s3_pipe_v;
		variable address: std_logic_vector(7 downto 0):="00000000";
		variable ro_addr_counter: integer range 0 to 131:=0;
		
		variable ro_flag: std_logic:='0';
		variable ram_counter: integer range 0 to 8:=0;
--		--========================================================		
		
	
	begin
		if rising_edge(clk_i) then
			if s3_pipeI.s2_pipe_data_mt22_o.s23_data_v_o='1' then
				s3_busy_o<='1';
				s3_pipe_wren_i<=x"F";
				s3_pipe_v.s3_pipe_mt22_data_v:=s3_pipeI.s2_pipe_data_mt22_o.s2_data_o;
				s3_pipe_v.s3_pipe_mt21_data_v:=s3_pipeI.s2_pipe_data_mt21_o.s2_data_o;
				s3_pipe_v.s3_pipe_mt12_data_v:=s3_pipeI.s2_pipe_data_mt12_o.s2_data_o;
				s3_pipe_v.s3_pipe_mt11_data_v:=s3_pipeI.s2_pipe_data_mt11_o.s2_data_o;
				
				s_data_port_arr_i(3)<=s3_pipe_v.s3_pipe_mt22_data_v;
				s_data_port_arr_i(2)<=s3_pipe_v.s3_pipe_mt21_data_v;
				s_data_port_arr_i(1)<=s3_pipe_v.s3_pipe_mt12_data_v;
				s_data_port_arr_i(0)<=s3_pipe_v.s3_pipe_mt11_data_v;
				
				if s3_flag < 128 then --Initiate s1 => s2 Readout
					if s3_flag=0 then
						s3_pipe_wren_i<=x"f";
						s3_flag := s3_flag +1; --increment counter
					
					else
						--Increment address ports of RAM modules
						s_addr_port_arr_i<= (others => (s_addr_port_arr_i(3) + 1));
						
						--Write new data to data ports of RAM modules

						s_data_port_arr_i(3)<=s3_pipe_v.s3_pipe_mt22_data_v;
						s_data_port_arr_i(2)<=s3_pipe_v.s3_pipe_mt21_data_v;
						s_data_port_arr_i(1)<=s3_pipe_v.s3_pipe_mt12_data_v;
						s_data_port_arr_i(0)<=s3_pipe_v.s3_pipe_mt11_data_v;
						
						--increment counter
						s3_flag := s3_flag +1; 
					end if;
				end if;
				
				elsif s3_flag = 128 then
					ro_flag:='1';
					s3_pipe_wren_i<=x"0";
					s_addr_port_arr_i<= (others =>"00000000");
				
				else -- if s2_flag=8 then --Flag end on s1 => s2 Readout
					s3_pipe_wren_i<=x"0";
					s_addr_port_arr_i<= (others =>"00000000");
				end if;
				--=================================================================
				if ro_flag='1' then
				case ram_counter is
					when 0 =>
						s3_pipe_rden_i<=x"1"; --Read enable on port a of ram 1
						s3_pipeO.s3_pipe_data_o<=s_data_port_arr_o(0); --Direct output data to sub ram data out
						case ro_addr_counter is 
							when 0 =>
								s_addr_port_arr_i(0)<=x"00";
								ro_addr_counter := ro_addr_counter + 1;
							when 1 =>
								s_addr_port_arr_i(0)<=x"01";
								ro_addr_counter := ro_addr_counter + 1;
							when 2 =>
								s_addr_port_arr_i(0)<=x"02";
								ro_addr_counter := ro_addr_counter + 1;
							when 3 =>
								s3_pipeO.s3_pipe_data_v_o<='1';
								s_addr_port_arr_i(0)<=x"03";
								ro_addr_counter := ro_addr_counter + 1;
							when 4 =>
								s_addr_port_arr_i(0)<=x"04";
								ro_addr_counter := ro_addr_counter + 1;
							when 5 =>
								s_addr_port_arr_i(0)<=x"05";
								ro_addr_counter := ro_addr_counter + 1;
							when 6 =>
								s_addr_port_arr_i(0)<=x"06";
								ro_addr_counter := ro_addr_counter + 1;
							when 7 =>
								s_addr_port_arr_i(0)<=x"07";
								ro_addr_counter := ro_addr_counter + 1;
							when 8 =>
								s_addr_port_arr_i(0)<=x"08";
								ro_addr_counter := ro_addr_counter + 1;
							when 9 =>
								s_addr_port_arr_i(0)<=x"09";
								ro_addr_counter := ro_addr_counter + 1;
							when 10 =>
								s_addr_port_arr_i(0)<=x"0A";
								ro_addr_counter := ro_addr_counter + 1;
							when 11 =>
								s_addr_port_arr_i(0)<=x"0B";
								ro_addr_counter := ro_addr_counter + 1;
							when 12 =>
								s_addr_port_arr_i(0)<=x"0C";
								ro_addr_counter := ro_addr_counter + 1;
							when 13 =>
								s_addr_port_arr_i(0)<=x"0D";
								ro_addr_counter := ro_addr_counter + 1;
							when 14 =>
								s_addr_port_arr_i(0)<=x"0E";
								ro_addr_counter := ro_addr_counter + 1;
							when 15 =>
								s_addr_port_arr_i(0)<=x"0F";
								ro_addr_counter := ro_addr_counter + 1;
							when 16 =>
								s_addr_port_arr_i(0)<=x"10";
								ro_addr_counter := ro_addr_counter + 1;
							when 17 =>
								s_addr_port_arr_i(0)<=x"11";
								ro_addr_counter := ro_addr_counter + 1;
							when 18 =>
								s_addr_port_arr_i(0)<=x"12";
								ro_addr_counter := ro_addr_counter + 1;
							when 19 =>
								s_addr_port_arr_i(0)<=x"13";
								ro_addr_counter := ro_addr_counter + 1;
							when 20 =>
								s_addr_port_arr_i(0)<=x"14";
								ro_addr_counter := ro_addr_counter + 1;
							when 21 =>
								s_addr_port_arr_i(0)<=x"15";
								ro_addr_counter := ro_addr_counter + 1;
							when 22 =>
								s_addr_port_arr_i(0)<=x"16";
								ro_addr_counter := ro_addr_counter + 1;
							when 23 =>
								s_addr_port_arr_i(0)<=x"17";
								ro_addr_counter := ro_addr_counter + 1;
							when 24 =>
								s_addr_port_arr_i(0)<=x"18";
								ro_addr_counter := ro_addr_counter + 1;
							when 25 =>
								s_addr_port_arr_i(0)<=x"19";
								ro_addr_counter := ro_addr_counter + 1;
							when 26 =>
								s_addr_port_arr_i(0)<=x"1A";
								ro_addr_counter := ro_addr_counter + 1;
							when 27 =>
								s_addr_port_arr_i(0)<=x"1B";
								ro_addr_counter := ro_addr_counter + 1;
							when 28 =>
								s_addr_port_arr_i(0)<=x"1C";
								ro_addr_counter := ro_addr_counter + 1;
							when 29 =>
								s_addr_port_arr_i(0)<=x"1D";
								ro_addr_counter := ro_addr_counter + 1;
							when 30 =>
								s_addr_port_arr_i(0)<=x"1E";
								ro_addr_counter := ro_addr_counter + 1;
							when 31 =>
								s_addr_port_arr_i(0)<=x"1F";
								ro_addr_counter := ro_addr_counter + 1;
							when 32 =>
								s_addr_port_arr_i(0)<=x"20";
								ro_addr_counter := ro_addr_counter + 1;
							when 33 =>
								s_addr_port_arr_i(0)<=x"21";
								ro_addr_counter := ro_addr_counter + 1;
							when 34 =>
								s_addr_port_arr_i(0)<=x"22";
								ro_addr_counter := ro_addr_counter + 1;
							when 35 =>
								s_addr_port_arr_i(0)<=x"23";
								ro_addr_counter := ro_addr_counter + 1;
							when 36 =>
								s_addr_port_arr_i(0)<=x"24";
								ro_addr_counter := ro_addr_counter + 1;
							when 37 =>
								s_addr_port_arr_i(0)<=x"25";
								ro_addr_counter := ro_addr_counter + 1;
							when 38 =>
								s_addr_port_arr_i(0)<=x"26";
								ro_addr_counter := ro_addr_counter + 1;
							when 39 =>
								s_addr_port_arr_i(0)<=x"27";
								ro_addr_counter := ro_addr_counter + 1;
							when 40 =>
								s_addr_port_arr_i(0)<=x"28";
								ro_addr_counter := ro_addr_counter + 1;
							when 41 =>
								s_addr_port_arr_i(0)<=x"29";
								ro_addr_counter := ro_addr_counter + 1;
							when 42 =>
								s_addr_port_arr_i(0)<=x"2A";
								ro_addr_counter := ro_addr_counter + 1;
							when 43 =>
								s_addr_port_arr_i(0)<=x"2B";
								ro_addr_counter := ro_addr_counter + 1;
							when 44 =>
								s_addr_port_arr_i(0)<=x"2C";
								ro_addr_counter := ro_addr_counter + 1;
							when 45 =>
								s_addr_port_arr_i(0)<=x"2D";
								ro_addr_counter := ro_addr_counter + 1;
							when 46 =>
								s_addr_port_arr_i(0)<=x"2E";
								ro_addr_counter := ro_addr_counter + 1;
							when 47 =>
								s_addr_port_arr_i(0)<=x"2F";
								ro_addr_counter := ro_addr_counter + 1;
							when 48 =>
								s_addr_port_arr_i(0)<=x"30";
								ro_addr_counter := ro_addr_counter + 1;
							when 49 =>
								s_addr_port_arr_i(0)<=x"31";
								ro_addr_counter := ro_addr_counter + 1;
							when 50 =>
								s_addr_port_arr_i(0)<=x"32";
								ro_addr_counter := ro_addr_counter + 1;
							when 51 =>
								s_addr_port_arr_i(0)<=x"33";
								ro_addr_counter := ro_addr_counter + 1;
							when 52 =>
								s_addr_port_arr_i(0)<=x"34";
								ro_addr_counter := ro_addr_counter + 1;
							when 53 =>
								s_addr_port_arr_i(0)<=x"35";
								ro_addr_counter := ro_addr_counter + 1;
							when 54 =>
								s_addr_port_arr_i(0)<=x"36";
								ro_addr_counter := ro_addr_counter + 1;
							when 55 =>
								s_addr_port_arr_i(0)<=x"37";
								ro_addr_counter := ro_addr_counter + 1;
							when 56 =>
								s_addr_port_arr_i(0)<=x"38";
								ro_addr_counter := ro_addr_counter + 1;
							when 57 =>
								s_addr_port_arr_i(0)<=x"39";
								ro_addr_counter := ro_addr_counter + 1;
							when 58 =>
								s_addr_port_arr_i(0)<=x"3A";
								ro_addr_counter := ro_addr_counter + 1;
							when 59 =>
								s_addr_port_arr_i(0)<=x"3B";
								ro_addr_counter := ro_addr_counter + 1;
							when 60 =>
								s_addr_port_arr_i(0)<=x"3C";
								ro_addr_counter := ro_addr_counter + 1;
							when 61 =>
								s_addr_port_arr_i(0)<=x"3D";
								ro_addr_counter := ro_addr_counter + 1;
							when 62 =>
								s_addr_port_arr_i(0)<=x"3E";
								ro_addr_counter := ro_addr_counter + 1;
							when 63 =>
								s_addr_port_arr_i(0)<=x"3F";
								ro_addr_counter := ro_addr_counter + 1;
							when 64 =>
								s_addr_port_arr_i(0)<=x"40";
								ro_addr_counter := ro_addr_counter + 1;
							when 65 =>
								s_addr_port_arr_i(0)<=x"41";
								ro_addr_counter := ro_addr_counter + 1;
							when 66 =>
								s_addr_port_arr_i(0)<=x"42";
								ro_addr_counter := ro_addr_counter + 1;
							when 67 =>
								s_addr_port_arr_i(0)<=x"43";
								ro_addr_counter := ro_addr_counter + 1;
							when 68 =>
								s_addr_port_arr_i(0)<=x"44";
								ro_addr_counter := ro_addr_counter + 1;
							when 69 =>
								s_addr_port_arr_i(0)<=x"45";
								ro_addr_counter := ro_addr_counter + 1;
							when 70 =>
								s_addr_port_arr_i(0)<=x"46";
								ro_addr_counter := ro_addr_counter + 1;
							when 71 =>
								s_addr_port_arr_i(0)<=x"47";
								ro_addr_counter := ro_addr_counter + 1;
							when 72 =>
								s_addr_port_arr_i(0)<=x"48";
								ro_addr_counter := ro_addr_counter + 1;
							when 73 =>
								s_addr_port_arr_i(0)<=x"49";
								ro_addr_counter := ro_addr_counter + 1;
							when 74 =>
								s_addr_port_arr_i(0)<=x"4A";
								ro_addr_counter := ro_addr_counter + 1;
							when 75 =>
								s_addr_port_arr_i(0)<=x"4B";
								ro_addr_counter := ro_addr_counter + 1;
							when 76 =>
								s_addr_port_arr_i(0)<=x"4C";
								ro_addr_counter := ro_addr_counter + 1;
							when 77 =>
								s_addr_port_arr_i(0)<=x"4D";
								ro_addr_counter := ro_addr_counter + 1;
							when 78 =>
								s_addr_port_arr_i(0)<=x"4E";
								ro_addr_counter := ro_addr_counter + 1;
							when 79 =>
								s_addr_port_arr_i(0)<=x"4F";
								ro_addr_counter := ro_addr_counter + 1;
							when 80 =>
								s_addr_port_arr_i(0)<=x"50";
								ro_addr_counter := ro_addr_counter + 1;
							when 81 =>
								s_addr_port_arr_i(0)<=x"51";
								ro_addr_counter := ro_addr_counter + 1;
							when 82 =>
								s_addr_port_arr_i(0)<=x"52";
								ro_addr_counter := ro_addr_counter + 1;
							when 83 =>
								s_addr_port_arr_i(0)<=x"53";
								ro_addr_counter := ro_addr_counter + 1;
							when 84 =>
								s_addr_port_arr_i(0)<=x"54";
								ro_addr_counter := ro_addr_counter + 1;
							when 85 =>
								s_addr_port_arr_i(0)<=x"55";
								ro_addr_counter := ro_addr_counter + 1;
							when 86 =>
								s_addr_port_arr_i(0)<=x"56";
								ro_addr_counter := ro_addr_counter + 1;
							when 87 =>
								s_addr_port_arr_i(0)<=x"57";
								ro_addr_counter := ro_addr_counter + 1;
							when 88 =>
								s_addr_port_arr_i(0)<=x"58";
								ro_addr_counter := ro_addr_counter + 1;
							when 89 =>
								s_addr_port_arr_i(0)<=x"59";
								ro_addr_counter := ro_addr_counter + 1;
							when 90 =>
								s_addr_port_arr_i(0)<=x"5A";
								ro_addr_counter := ro_addr_counter + 1;
							when 91 =>
								s_addr_port_arr_i(0)<=x"5B";
								ro_addr_counter := ro_addr_counter + 1;
							when 92 =>
								s_addr_port_arr_i(0)<=x"5C";
								ro_addr_counter := ro_addr_counter + 1;
							when 93 =>
								s_addr_port_arr_i(0)<=x"5D";
								ro_addr_counter := ro_addr_counter + 1;
							when 94 =>
								s_addr_port_arr_i(0)<=x"5E";
								ro_addr_counter := ro_addr_counter + 1;
							when 95 =>
								s_addr_port_arr_i(0)<=x"5F";
								ro_addr_counter := ro_addr_counter + 1;
							when 96 =>
								s_addr_port_arr_i(0)<=x"60";
								ro_addr_counter := ro_addr_counter + 1;
							when 97 =>
								s_addr_port_arr_i(0)<=x"61";
								ro_addr_counter := ro_addr_counter + 1;
							when 98 =>
								s_addr_port_arr_i(0)<=x"62";
								ro_addr_counter := ro_addr_counter + 1;
							when 99 =>
								s_addr_port_arr_i(0)<=x"63";
								ro_addr_counter := ro_addr_counter + 1;
							when 100 =>
								s_addr_port_arr_i(0)<=x"64";
								ro_addr_counter := ro_addr_counter + 1;
							when 101 =>
								s_addr_port_arr_i(0)<=x"65";
								ro_addr_counter := ro_addr_counter + 1;
							when 102 =>
								s_addr_port_arr_i(0)<=x"66";
								ro_addr_counter := ro_addr_counter + 1;
							when 103 =>
								s_addr_port_arr_i(0)<=x"67";
								ro_addr_counter := ro_addr_counter + 1;
							when 104 =>
								s_addr_port_arr_i(0)<=x"68";
								ro_addr_counter := ro_addr_counter + 1;
							when 105 =>
								s_addr_port_arr_i(0)<=x"69";
								ro_addr_counter := ro_addr_counter + 1;
							when 106 =>
								s_addr_port_arr_i(0)<=x"6A";
								ro_addr_counter := ro_addr_counter + 1;
							when 107 =>
								s_addr_port_arr_i(0)<=x"6B";
								ro_addr_counter := ro_addr_counter + 1;
							when 108 =>
								s_addr_port_arr_i(0)<=x"6C";
								ro_addr_counter := ro_addr_counter + 1;
							when 109 =>
								s_addr_port_arr_i(0)<=x"6D";
								ro_addr_counter := ro_addr_counter + 1;
							when 110 =>
								s_addr_port_arr_i(0)<=x"6E";
								ro_addr_counter := ro_addr_counter + 1;
							when 111 =>
								s_addr_port_arr_i(0)<=x"6F";
								ro_addr_counter := ro_addr_counter + 1;
							when 112 =>
								s_addr_port_arr_i(0)<=x"70";
								ro_addr_counter := ro_addr_counter + 1;
							when 113 =>
								s_addr_port_arr_i(0)<=x"71";
								ro_addr_counter := ro_addr_counter + 1;
							when 114 =>
								s_addr_port_arr_i(0)<=x"72";
								ro_addr_counter := ro_addr_counter + 1;
							when 115 =>
								s_addr_port_arr_i(0)<=x"73";
								ro_addr_counter := ro_addr_counter + 1;
							when 116 =>
								s_addr_port_arr_i(0)<=x"74";
								ro_addr_counter := ro_addr_counter + 1;
							when 117 =>
								s_addr_port_arr_i(0)<=x"75";
								ro_addr_counter := ro_addr_counter + 1;
							when 118 =>
								s_addr_port_arr_i(0)<=x"76";
								ro_addr_counter := ro_addr_counter + 1;
							when 119 =>
								s_addr_port_arr_i(0)<=x"77";
								ro_addr_counter := ro_addr_counter + 1;
							when 120 =>
								s_addr_port_arr_i(0)<=x"78";
								ro_addr_counter := ro_addr_counter + 1;
							when 121 =>
								s_addr_port_arr_i(0)<=x"79";
								ro_addr_counter := ro_addr_counter + 1;
							when 122 =>
								s_addr_port_arr_i(0)<=x"7A";
								ro_addr_counter := ro_addr_counter + 1;
							when 123 =>
								s_addr_port_arr_i(0)<=x"7B";
								ro_addr_counter := ro_addr_counter + 1;
							when 124 =>
								s_addr_port_arr_i(0)<=x"7C";
								ro_addr_counter := ro_addr_counter + 1;
							when 125 =>
								s_addr_port_arr_i(0)<=x"7D";
								ro_addr_counter := ro_addr_counter + 1;
							when 126 =>
								s_addr_port_arr_i(0)<=x"7E";
								ro_addr_counter := ro_addr_counter + 1;
							when 127 =>
								s_addr_port_arr_i(0)<=x"7F";
								ro_addr_counter := ro_addr_counter + 1;
							when 128 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"2"; --Read enable on port a of ram 2
								s_addr_port_arr_i(1)<=x"00";
							when 129 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"2"; --Read enable on port a of ram 2
								s_addr_port_arr_i(1)<=x"01";
							when 130 =>
								ro_addr_counter := 0;
								s3_pipe_rden_i<=x"2"; --Read enable on port a of ram 2
								s_addr_port_arr_i(1)<=x"02";
								ram_counter:= ram_counter + 1; --Increment RAM counter
							when others =>
						end case;
					when 1 =>
						s3_pipe_rden_i<=x"2"; --Read enable on port a of ram 2
						s3_pipeO.s3_pipe_data_o<=s_data_port_arr_o(1); --Direct output data to sub ram data out
						case ro_addr_counter is 
							when 0 =>
								s_addr_port_arr_i(1)<=x"03";
								ro_addr_counter := ro_addr_counter + 1;
							when 1 =>
								s_addr_port_arr_i(1)<=x"04";
								ro_addr_counter := ro_addr_counter + 1;
							when 2 =>
								s_addr_port_arr_i(1)<=x"05";
								ro_addr_counter := ro_addr_counter + 1;
							when 3 =>
								s_addr_port_arr_i(1)<=x"06";
								ro_addr_counter := ro_addr_counter + 1;
							when 4 =>
								s_addr_port_arr_i(1)<=x"07";
								ro_addr_counter := ro_addr_counter + 1;
							when 5 =>
								s_addr_port_arr_i(1)<=x"08";
								ro_addr_counter := ro_addr_counter + 1;
							when 6 =>
								s_addr_port_arr_i(1)<=x"09";
								ro_addr_counter := ro_addr_counter + 1;
							when 7 =>
								s_addr_port_arr_i(1)<=x"0A";
								ro_addr_counter := ro_addr_counter + 1;
							when 8 =>
								s_addr_port_arr_i(1)<=x"0B";
								ro_addr_counter := ro_addr_counter + 1;
							when 9 =>
								s_addr_port_arr_i(1)<=x"0C";
								ro_addr_counter := ro_addr_counter + 1;
							when 10 =>
								s_addr_port_arr_i(1)<=x"0D";
								ro_addr_counter := ro_addr_counter + 1;
							when 11 =>
								s_addr_port_arr_i(1)<=x"0E";
								ro_addr_counter := ro_addr_counter + 1;
							when 12 =>
								s_addr_port_arr_i(1)<=x"0F";
								ro_addr_counter := ro_addr_counter + 1;
							when 13 =>
								s_addr_port_arr_i(1)<=x"10";
								ro_addr_counter := ro_addr_counter + 1;
							when 14 =>
								s_addr_port_arr_i(1)<=x"11";
								ro_addr_counter := ro_addr_counter + 1;
							when 15 =>
								s_addr_port_arr_i(1)<=x"12";
								ro_addr_counter := ro_addr_counter + 1;
							when 16 =>
								s_addr_port_arr_i(1)<=x"13";
								ro_addr_counter := ro_addr_counter + 1;
							when 17 =>
								s_addr_port_arr_i(1)<=x"14";
								ro_addr_counter := ro_addr_counter + 1;
							when 18 =>
								s_addr_port_arr_i(1)<=x"15";
								ro_addr_counter := ro_addr_counter + 1;
							when 19 =>
								s_addr_port_arr_i(1)<=x"16";
								ro_addr_counter := ro_addr_counter + 1;
							when 20 =>
								s_addr_port_arr_i(1)<=x"17";
								ro_addr_counter := ro_addr_counter + 1;
							when 21 =>
								s_addr_port_arr_i(1)<=x"18";
								ro_addr_counter := ro_addr_counter + 1;
							when 22 =>
								s_addr_port_arr_i(1)<=x"19";
								ro_addr_counter := ro_addr_counter + 1;
							when 23 =>
								s_addr_port_arr_i(1)<=x"1A";
								ro_addr_counter := ro_addr_counter + 1;
							when 24 =>
								s_addr_port_arr_i(1)<=x"1B";
								ro_addr_counter := ro_addr_counter + 1;
							when 25 =>
								s_addr_port_arr_i(1)<=x"1C";
								ro_addr_counter := ro_addr_counter + 1;
							when 26 =>
								s_addr_port_arr_i(1)<=x"1D";
								ro_addr_counter := ro_addr_counter + 1;
							when 27 =>
								s_addr_port_arr_i(1)<=x"1E";
								ro_addr_counter := ro_addr_counter + 1;
							when 28 =>
								s_addr_port_arr_i(1)<=x"1F";
								ro_addr_counter := ro_addr_counter + 1;
							when 29 =>
								s_addr_port_arr_i(1)<=x"20";
								ro_addr_counter := ro_addr_counter + 1;
							when 30 =>
								s_addr_port_arr_i(1)<=x"21";
								ro_addr_counter := ro_addr_counter + 1;
							when 31 =>
								s_addr_port_arr_i(1)<=x"22";
								ro_addr_counter := ro_addr_counter + 1;
							when 32 =>
								s_addr_port_arr_i(1)<=x"23";
								ro_addr_counter := ro_addr_counter + 1;
							when 33 =>
								s_addr_port_arr_i(1)<=x"24";
								ro_addr_counter := ro_addr_counter + 1;
							when 34 =>
								s_addr_port_arr_i(1)<=x"25";
								ro_addr_counter := ro_addr_counter + 1;
							when 35 =>
								s_addr_port_arr_i(1)<=x"26";
								ro_addr_counter := ro_addr_counter + 1;
							when 36 =>
								s_addr_port_arr_i(1)<=x"27";
								ro_addr_counter := ro_addr_counter + 1;
							when 37 =>
								s_addr_port_arr_i(1)<=x"28";
								ro_addr_counter := ro_addr_counter + 1;
							when 38 =>
								s_addr_port_arr_i(1)<=x"29";
								ro_addr_counter := ro_addr_counter + 1;
							when 39 =>
								s_addr_port_arr_i(1)<=x"2A";
								ro_addr_counter := ro_addr_counter + 1;
							when 40 =>
								s_addr_port_arr_i(1)<=x"2B";
								ro_addr_counter := ro_addr_counter + 1;
							when 41 =>
								s_addr_port_arr_i(1)<=x"2C";
								ro_addr_counter := ro_addr_counter + 1;
							when 42 =>
								s_addr_port_arr_i(1)<=x"2D";
								ro_addr_counter := ro_addr_counter + 1;
							when 43 =>
								s_addr_port_arr_i(1)<=x"2E";
								ro_addr_counter := ro_addr_counter + 1;
							when 44 =>
								s_addr_port_arr_i(1)<=x"2F";
								ro_addr_counter := ro_addr_counter + 1;
							when 45 =>
								s_addr_port_arr_i(1)<=x"30";
								ro_addr_counter := ro_addr_counter + 1;
							when 46 =>
								s_addr_port_arr_i(1)<=x"31";
								ro_addr_counter := ro_addr_counter + 1;
							when 47 =>
								s_addr_port_arr_i(1)<=x"32";
								ro_addr_counter := ro_addr_counter + 1;
							when 48 =>
								s_addr_port_arr_i(1)<=x"33";
								ro_addr_counter := ro_addr_counter + 1;
							when 49 =>
								s_addr_port_arr_i(1)<=x"34";
								ro_addr_counter := ro_addr_counter + 1;
							when 50 =>
								s_addr_port_arr_i(1)<=x"35";
								ro_addr_counter := ro_addr_counter + 1;
							when 51 =>
								s_addr_port_arr_i(1)<=x"36";
								ro_addr_counter := ro_addr_counter + 1;
							when 52 =>
								s_addr_port_arr_i(1)<=x"37";
								ro_addr_counter := ro_addr_counter + 1;
							when 53 =>
								s_addr_port_arr_i(1)<=x"38";
								ro_addr_counter := ro_addr_counter + 1;
							when 54 =>
								s_addr_port_arr_i(1)<=x"39";
								ro_addr_counter := ro_addr_counter + 1;
							when 55 =>
								s_addr_port_arr_i(1)<=x"3A";
								ro_addr_counter := ro_addr_counter + 1;
							when 56 =>
								s_addr_port_arr_i(1)<=x"3B";
								ro_addr_counter := ro_addr_counter + 1;
							when 57 =>
								s_addr_port_arr_i(1)<=x"3C";
								ro_addr_counter := ro_addr_counter + 1;
							when 58 =>
								s_addr_port_arr_i(1)<=x"3D";
								ro_addr_counter := ro_addr_counter + 1;
							when 59 =>
								s_addr_port_arr_i(1)<=x"3E";
								ro_addr_counter := ro_addr_counter + 1;
							when 60 =>
								s_addr_port_arr_i(1)<=x"3F";
								ro_addr_counter := ro_addr_counter + 1;
							when 61 =>
								s_addr_port_arr_i(1)<=x"40";
								ro_addr_counter := ro_addr_counter + 1;
							when 62 =>
								s_addr_port_arr_i(1)<=x"41";
								ro_addr_counter := ro_addr_counter + 1;
							when 63 =>
								s_addr_port_arr_i(1)<=x"42";
								ro_addr_counter := ro_addr_counter + 1;
							when 64 =>
								s_addr_port_arr_i(1)<=x"43";
								ro_addr_counter := ro_addr_counter + 1;
							when 65 =>
								s_addr_port_arr_i(1)<=x"44";
								ro_addr_counter := ro_addr_counter + 1;
							when 66 =>
								s_addr_port_arr_i(1)<=x"45";
								ro_addr_counter := ro_addr_counter + 1;
							when 67 =>
								s_addr_port_arr_i(1)<=x"46";
								ro_addr_counter := ro_addr_counter + 1;
							when 68 =>
								s_addr_port_arr_i(1)<=x"47";
								ro_addr_counter := ro_addr_counter + 1;
							when 69 =>
								s_addr_port_arr_i(1)<=x"48";
								ro_addr_counter := ro_addr_counter + 1;
							when 70 =>
								s_addr_port_arr_i(1)<=x"49";
								ro_addr_counter := ro_addr_counter + 1;
							when 71 =>
								s_addr_port_arr_i(1)<=x"4A";
								ro_addr_counter := ro_addr_counter + 1;
							when 72 =>
								s_addr_port_arr_i(1)<=x"4B";
								ro_addr_counter := ro_addr_counter + 1;
							when 73 =>
								s_addr_port_arr_i(1)<=x"4C";
								ro_addr_counter := ro_addr_counter + 1;
							when 74 =>
								s_addr_port_arr_i(1)<=x"4D";
								ro_addr_counter := ro_addr_counter + 1;
							when 75 =>
								s_addr_port_arr_i(1)<=x"4E";
								ro_addr_counter := ro_addr_counter + 1;
							when 76 =>
								s_addr_port_arr_i(1)<=x"4F";
								ro_addr_counter := ro_addr_counter + 1;
							when 77 =>
								s_addr_port_arr_i(1)<=x"50";
								ro_addr_counter := ro_addr_counter + 1;
							when 78 =>
								s_addr_port_arr_i(1)<=x"51";
								ro_addr_counter := ro_addr_counter + 1;
							when 79 =>
								s_addr_port_arr_i(1)<=x"52";
								ro_addr_counter := ro_addr_counter + 1;
							when 80 =>
								s_addr_port_arr_i(1)<=x"53";
								ro_addr_counter := ro_addr_counter + 1;
							when 81 =>
								s_addr_port_arr_i(1)<=x"54";
								ro_addr_counter := ro_addr_counter + 1;
							when 82 =>
								s_addr_port_arr_i(1)<=x"55";
								ro_addr_counter := ro_addr_counter + 1;
							when 83 =>
								s_addr_port_arr_i(1)<=x"56";
								ro_addr_counter := ro_addr_counter + 1;
							when 84 =>
								s_addr_port_arr_i(1)<=x"57";
								ro_addr_counter := ro_addr_counter + 1;
							when 85 =>
								s_addr_port_arr_i(1)<=x"58";
								ro_addr_counter := ro_addr_counter + 1;
							when 86 =>
								s_addr_port_arr_i(1)<=x"59";
								ro_addr_counter := ro_addr_counter + 1;
							when 87 =>
								s_addr_port_arr_i(1)<=x"5A";
								ro_addr_counter := ro_addr_counter + 1;
							when 88 =>
								s_addr_port_arr_i(1)<=x"5B";
								ro_addr_counter := ro_addr_counter + 1;
							when 89 =>
								s_addr_port_arr_i(1)<=x"5C";
								ro_addr_counter := ro_addr_counter + 1;
							when 90 =>
								s_addr_port_arr_i(1)<=x"5D";
								ro_addr_counter := ro_addr_counter + 1;
							when 91 =>
								s_addr_port_arr_i(1)<=x"5E";
								ro_addr_counter := ro_addr_counter + 1;
							when 92 =>
								s_addr_port_arr_i(1)<=x"5F";
								ro_addr_counter := ro_addr_counter + 1;
							when 93 =>
								s_addr_port_arr_i(1)<=x"60";
								ro_addr_counter := ro_addr_counter + 1;
							when 94 =>
								s_addr_port_arr_i(1)<=x"61";
								ro_addr_counter := ro_addr_counter + 1;
							when 95 =>
								s_addr_port_arr_i(1)<=x"62";
								ro_addr_counter := ro_addr_counter + 1;
							when 96 =>
								s_addr_port_arr_i(1)<=x"63";
								ro_addr_counter := ro_addr_counter + 1;
							when 97 =>
								s_addr_port_arr_i(1)<=x"64";
								ro_addr_counter := ro_addr_counter + 1;
							when 98 =>
								s_addr_port_arr_i(1)<=x"65";
								ro_addr_counter := ro_addr_counter + 1;
							when 99 =>
								s_addr_port_arr_i(1)<=x"66";
								ro_addr_counter := ro_addr_counter + 1;
							when 100 =>
								s_addr_port_arr_i(1)<=x"67";
								ro_addr_counter := ro_addr_counter + 1;
							when 101 =>
								s_addr_port_arr_i(1)<=x"68";
								ro_addr_counter := ro_addr_counter + 1;
							when 102 =>
								s_addr_port_arr_i(1)<=x"69";
								ro_addr_counter := ro_addr_counter + 1;
							when 103 =>
								s_addr_port_arr_i(1)<=x"6A";
								ro_addr_counter := ro_addr_counter + 1;
							when 104 =>
								s_addr_port_arr_i(1)<=x"6B";
								ro_addr_counter := ro_addr_counter + 1;
							when 105 =>
								s_addr_port_arr_i(1)<=x"6C";
								ro_addr_counter := ro_addr_counter + 1;
							when 106 =>
								s_addr_port_arr_i(1)<=x"6D";
								ro_addr_counter := ro_addr_counter + 1;
							when 107 =>
								s_addr_port_arr_i(1)<=x"6E";
								ro_addr_counter := ro_addr_counter + 1;
							when 108 =>
								s_addr_port_arr_i(1)<=x"6F";
								ro_addr_counter := ro_addr_counter + 1;
							when 109 =>
								s_addr_port_arr_i(1)<=x"70";
								ro_addr_counter := ro_addr_counter + 1;
							when 110 =>
								s_addr_port_arr_i(1)<=x"71";
								ro_addr_counter := ro_addr_counter + 1;
							when 111 =>
								s_addr_port_arr_i(1)<=x"72";
								ro_addr_counter := ro_addr_counter + 1;
							when 112 =>
								s_addr_port_arr_i(1)<=x"73";
								ro_addr_counter := ro_addr_counter + 1;
							when 113 =>
								s_addr_port_arr_i(1)<=x"74";
								ro_addr_counter := ro_addr_counter + 1;
							when 114 =>
								s_addr_port_arr_i(1)<=x"75";
								ro_addr_counter := ro_addr_counter + 1;
							when 115 =>
								s_addr_port_arr_i(1)<=x"76";
								ro_addr_counter := ro_addr_counter + 1;
							when 116 =>
								s_addr_port_arr_i(1)<=x"77";
								ro_addr_counter := ro_addr_counter + 1;
							when 117 =>
								s_addr_port_arr_i(1)<=x"78";
								ro_addr_counter := ro_addr_counter + 1;
							when 118 =>
								s_addr_port_arr_i(1)<=x"79";
								ro_addr_counter := ro_addr_counter + 1;
							when 119 =>
								s_addr_port_arr_i(1)<=x"7A";
								ro_addr_counter := ro_addr_counter + 1;
							when 120 =>
								s_addr_port_arr_i(1)<=x"7B";
								ro_addr_counter := ro_addr_counter + 1;
							when 121 =>
								s_addr_port_arr_i(1)<=x"7C";
								ro_addr_counter := ro_addr_counter + 1;
							when 122 =>
								s_addr_port_arr_i(1)<=x"7D";
								ro_addr_counter := ro_addr_counter + 1;
							when 123 =>
								s_addr_port_arr_i(1)<=x"7E";
								ro_addr_counter := ro_addr_counter + 1;
							when 124 =>
								s_addr_port_arr_i(1)<=x"7F";
								ro_addr_counter := ro_addr_counter + 1;
							when 125 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"4"; --Read enable on port a of ram 2
								s_addr_port_arr_i(2)<=x"00";
							when 126 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"4"; --Read enable on port a of ram 2
								s_addr_port_arr_i(2)<=x"01";
							when 127 =>
							ro_addr_counter := 0;
								s3_pipe_rden_i<=x"4";--Read enable on port a of ram 2
								s_addr_port_arr_i(2)<=x"02";
								ram_counter:= ram_counter + 1; --Increment RAM counter
							when others =>
						end case;
					when 2 =>
						s3_pipe_rden_i<=x"4"; --Read enable on port a of ram 3
						s3_pipeO.s3_pipe_data_o<=s_data_port_arr_o(2); --Direct output data to sub ram data out
						case ro_addr_counter is 
							when 0 =>
								s_addr_port_arr_i(2)<=x"03";
								ro_addr_counter := ro_addr_counter + 1;
							when 1 =>
								s_addr_port_arr_i(2)<=x"04";
								ro_addr_counter := ro_addr_counter + 1;
							when 2 =>
								s_addr_port_arr_i(2)<=x"05";
								ro_addr_counter := ro_addr_counter + 1;
							when 3 =>
								s_addr_port_arr_i(2)<=x"06";
								ro_addr_counter := ro_addr_counter + 1;
							when 4 =>
								s_addr_port_arr_i(2)<=x"07";
								ro_addr_counter := ro_addr_counter + 1;
							when 5 =>
								s_addr_port_arr_i(2)<=x"08";
								ro_addr_counter := ro_addr_counter + 1;
							when 6 =>
								s_addr_port_arr_i(2)<=x"09";
								ro_addr_counter := ro_addr_counter + 1;
							when 7 =>
								s_addr_port_arr_i(2)<=x"0A";
								ro_addr_counter := ro_addr_counter + 1;
							when 8 =>
								s_addr_port_arr_i(2)<=x"0B";
								ro_addr_counter := ro_addr_counter + 1;
							when 9 =>
								s_addr_port_arr_i(2)<=x"0C";
								ro_addr_counter := ro_addr_counter + 1;
							when 10 =>
								s_addr_port_arr_i(2)<=x"0D";
								ro_addr_counter := ro_addr_counter + 1;
							when 11 =>
								s_addr_port_arr_i(2)<=x"0E";
								ro_addr_counter := ro_addr_counter + 1;
							when 12 =>
								s_addr_port_arr_i(2)<=x"0F";
								ro_addr_counter := ro_addr_counter + 1;
							when 13 =>
								s_addr_port_arr_i(2)<=x"10";
								ro_addr_counter := ro_addr_counter + 1;
							when 14 =>
								s_addr_port_arr_i(2)<=x"11";
								ro_addr_counter := ro_addr_counter + 1;
							when 15 =>
								s_addr_port_arr_i(2)<=x"12";
								ro_addr_counter := ro_addr_counter + 1;
							when 16 =>
								s_addr_port_arr_i(2)<=x"13";
								ro_addr_counter := ro_addr_counter + 1;
							when 17 =>
								s_addr_port_arr_i(2)<=x"14";
								ro_addr_counter := ro_addr_counter + 1;
							when 18 =>
								s_addr_port_arr_i(2)<=x"15";
								ro_addr_counter := ro_addr_counter + 1;
							when 19 =>
								s_addr_port_arr_i(2)<=x"16";
								ro_addr_counter := ro_addr_counter + 1;
							when 20 =>
								s_addr_port_arr_i(2)<=x"17";
								ro_addr_counter := ro_addr_counter + 1;
							when 21 =>
								s_addr_port_arr_i(2)<=x"18";
								ro_addr_counter := ro_addr_counter + 1;
							when 22 =>
								s_addr_port_arr_i(2)<=x"19";
								ro_addr_counter := ro_addr_counter + 1;
							when 23 =>
								s_addr_port_arr_i(2)<=x"1A";
								ro_addr_counter := ro_addr_counter + 1;
							when 24 =>
								s_addr_port_arr_i(2)<=x"1B";
								ro_addr_counter := ro_addr_counter + 1;
							when 25 =>
								s_addr_port_arr_i(2)<=x"1C";
								ro_addr_counter := ro_addr_counter + 1;
							when 26 =>
								s_addr_port_arr_i(2)<=x"1D";
								ro_addr_counter := ro_addr_counter + 1;
							when 27 =>
								s_addr_port_arr_i(2)<=x"1E";
								ro_addr_counter := ro_addr_counter + 1;
							when 28 =>
								s_addr_port_arr_i(2)<=x"1F";
								ro_addr_counter := ro_addr_counter + 1;
							when 29 =>
								s_addr_port_arr_i(2)<=x"20";
								ro_addr_counter := ro_addr_counter + 1;
							when 30 =>
								s_addr_port_arr_i(2)<=x"21";
								ro_addr_counter := ro_addr_counter + 1;
							when 31 =>
								s_addr_port_arr_i(2)<=x"22";
								ro_addr_counter := ro_addr_counter + 1;
							when 32 =>
								s_addr_port_arr_i(2)<=x"23";
								ro_addr_counter := ro_addr_counter + 1;
							when 33 =>
								s_addr_port_arr_i(2)<=x"24";
								ro_addr_counter := ro_addr_counter + 1;
							when 34 =>
								s_addr_port_arr_i(2)<=x"25";
								ro_addr_counter := ro_addr_counter + 1;
							when 35 =>
								s_addr_port_arr_i(2)<=x"26";
								ro_addr_counter := ro_addr_counter + 1;
							when 36 =>
								s_addr_port_arr_i(2)<=x"27";
								ro_addr_counter := ro_addr_counter + 1;
							when 37 =>
								s_addr_port_arr_i(2)<=x"28";
								ro_addr_counter := ro_addr_counter + 1;
							when 38 =>
								s_addr_port_arr_i(2)<=x"29";
								ro_addr_counter := ro_addr_counter + 1;
							when 39 =>
								s_addr_port_arr_i(2)<=x"2A";
								ro_addr_counter := ro_addr_counter + 1;
							when 40 =>
								s_addr_port_arr_i(2)<=x"2B";
								ro_addr_counter := ro_addr_counter + 1;
							when 41 =>
								s_addr_port_arr_i(2)<=x"2C";
								ro_addr_counter := ro_addr_counter + 1;
							when 42 =>
								s_addr_port_arr_i(2)<=x"2D";
								ro_addr_counter := ro_addr_counter + 1;
							when 43 =>
								s_addr_port_arr_i(2)<=x"2E";
								ro_addr_counter := ro_addr_counter + 1;
							when 44 =>
								s_addr_port_arr_i(2)<=x"2F";
								ro_addr_counter := ro_addr_counter + 1;
							when 45 =>
								s_addr_port_arr_i(2)<=x"30";
								ro_addr_counter := ro_addr_counter + 1;
							when 46 =>
								s_addr_port_arr_i(2)<=x"31";
								ro_addr_counter := ro_addr_counter + 1;
							when 47 =>
								s_addr_port_arr_i(2)<=x"32";
								ro_addr_counter := ro_addr_counter + 1;
							when 48 =>
								s_addr_port_arr_i(2)<=x"33";
								ro_addr_counter := ro_addr_counter + 1;
							when 49 =>
								s_addr_port_arr_i(2)<=x"34";
								ro_addr_counter := ro_addr_counter + 1;
							when 50 =>
								s_addr_port_arr_i(2)<=x"35";
								ro_addr_counter := ro_addr_counter + 1;
							when 51 =>
								s_addr_port_arr_i(2)<=x"36";
								ro_addr_counter := ro_addr_counter + 1;
							when 52 =>
								s_addr_port_arr_i(2)<=x"37";
								ro_addr_counter := ro_addr_counter + 1;
							when 53 =>
								s_addr_port_arr_i(2)<=x"38";
								ro_addr_counter := ro_addr_counter + 1;
							when 54 =>
								s_addr_port_arr_i(2)<=x"39";
								ro_addr_counter := ro_addr_counter + 1;
							when 55 =>
								s_addr_port_arr_i(2)<=x"3A";
								ro_addr_counter := ro_addr_counter + 1;
							when 56 =>
								s_addr_port_arr_i(2)<=x"3B";
								ro_addr_counter := ro_addr_counter + 1;
							when 57 =>
								s_addr_port_arr_i(2)<=x"3C";
								ro_addr_counter := ro_addr_counter + 1;
							when 58 =>
								s_addr_port_arr_i(2)<=x"3D";
								ro_addr_counter := ro_addr_counter + 1;
							when 59 =>
								s_addr_port_arr_i(2)<=x"3E";
								ro_addr_counter := ro_addr_counter + 1;
							when 60 =>
								s_addr_port_arr_i(2)<=x"3F";
								ro_addr_counter := ro_addr_counter + 1;
							when 61 =>
								s_addr_port_arr_i(2)<=x"40";
								ro_addr_counter := ro_addr_counter + 1;
							when 62 =>
								s_addr_port_arr_i(2)<=x"41";
								ro_addr_counter := ro_addr_counter + 1;
							when 63 =>
								s_addr_port_arr_i(2)<=x"42";
								ro_addr_counter := ro_addr_counter + 1;
							when 64 =>
								s_addr_port_arr_i(2)<=x"43";
								ro_addr_counter := ro_addr_counter + 1;
							when 65 =>
								s_addr_port_arr_i(2)<=x"44";
								ro_addr_counter := ro_addr_counter + 1;
							when 66 =>
								s_addr_port_arr_i(2)<=x"45";
								ro_addr_counter := ro_addr_counter + 1;
							when 67 =>
								s_addr_port_arr_i(2)<=x"46";
								ro_addr_counter := ro_addr_counter + 1;
							when 68 =>
								s_addr_port_arr_i(2)<=x"47";
								ro_addr_counter := ro_addr_counter + 1;
							when 69 =>
								s_addr_port_arr_i(2)<=x"48";
								ro_addr_counter := ro_addr_counter + 1;
							when 70 =>
								s_addr_port_arr_i(2)<=x"49";
								ro_addr_counter := ro_addr_counter + 1;
							when 71 =>
								s_addr_port_arr_i(2)<=x"4A";
								ro_addr_counter := ro_addr_counter + 1;
							when 72 =>
								s_addr_port_arr_i(2)<=x"4B";
								ro_addr_counter := ro_addr_counter + 1;
							when 73 =>
								s_addr_port_arr_i(2)<=x"4C";
								ro_addr_counter := ro_addr_counter + 1;
							when 74 =>
								s_addr_port_arr_i(2)<=x"4D";
								ro_addr_counter := ro_addr_counter + 1;
							when 75 =>
								s_addr_port_arr_i(2)<=x"4E";
								ro_addr_counter := ro_addr_counter + 1;
							when 76 =>
								s_addr_port_arr_i(2)<=x"4F";
								ro_addr_counter := ro_addr_counter + 1;
							when 77 =>
								s_addr_port_arr_i(2)<=x"50";
								ro_addr_counter := ro_addr_counter + 1;
							when 78 =>
								s_addr_port_arr_i(2)<=x"51";
								ro_addr_counter := ro_addr_counter + 1;
							when 79 =>
								s_addr_port_arr_i(2)<=x"52";
								ro_addr_counter := ro_addr_counter + 1;
							when 80 =>
								s_addr_port_arr_i(2)<=x"53";
								ro_addr_counter := ro_addr_counter + 1;
							when 81 =>
								s_addr_port_arr_i(2)<=x"54";
								ro_addr_counter := ro_addr_counter + 1;
							when 82 =>
								s_addr_port_arr_i(2)<=x"55";
								ro_addr_counter := ro_addr_counter + 1;
							when 83 =>
								s_addr_port_arr_i(2)<=x"56";
								ro_addr_counter := ro_addr_counter + 1;
							when 84 =>
								s_addr_port_arr_i(2)<=x"57";
								ro_addr_counter := ro_addr_counter + 1;
							when 85 =>
								s_addr_port_arr_i(2)<=x"58";
								ro_addr_counter := ro_addr_counter + 1;
							when 86 =>
								s_addr_port_arr_i(2)<=x"59";
								ro_addr_counter := ro_addr_counter + 1;
							when 87 =>
								s_addr_port_arr_i(2)<=x"5A";
								ro_addr_counter := ro_addr_counter + 1;
							when 88 =>
								s_addr_port_arr_i(2)<=x"5B";
								ro_addr_counter := ro_addr_counter + 1;
							when 89 =>
								s_addr_port_arr_i(2)<=x"5C";
								ro_addr_counter := ro_addr_counter + 1;
							when 90 =>
								s_addr_port_arr_i(2)<=x"5D";
								ro_addr_counter := ro_addr_counter + 1;
							when 91 =>
								s_addr_port_arr_i(2)<=x"5E";
								ro_addr_counter := ro_addr_counter + 1;
							when 92 =>
								s_addr_port_arr_i(2)<=x"5F";
								ro_addr_counter := ro_addr_counter + 1;
							when 93 =>
								s_addr_port_arr_i(2)<=x"60";
								ro_addr_counter := ro_addr_counter + 1;
							when 94 =>
								s_addr_port_arr_i(2)<=x"61";
								ro_addr_counter := ro_addr_counter + 1;
							when 95 =>
								s_addr_port_arr_i(2)<=x"62";
								ro_addr_counter := ro_addr_counter + 1;
							when 96 =>
								s_addr_port_arr_i(2)<=x"63";
								ro_addr_counter := ro_addr_counter + 1;
							when 97 =>
								s_addr_port_arr_i(2)<=x"64";
								ro_addr_counter := ro_addr_counter + 1;
							when 98 =>
								s_addr_port_arr_i(2)<=x"65";
								ro_addr_counter := ro_addr_counter + 1;
							when 99 =>
								s_addr_port_arr_i(2)<=x"66";
								ro_addr_counter := ro_addr_counter + 1;
							when 100 =>
								s_addr_port_arr_i(2)<=x"67";
								ro_addr_counter := ro_addr_counter + 1;
							when 101 =>
								s_addr_port_arr_i(2)<=x"68";
								ro_addr_counter := ro_addr_counter + 1;
							when 102 =>
								s_addr_port_arr_i(2)<=x"69";
								ro_addr_counter := ro_addr_counter + 1;
							when 103 =>
								s_addr_port_arr_i(2)<=x"6A";
								ro_addr_counter := ro_addr_counter + 1;
							when 104 =>
								s_addr_port_arr_i(2)<=x"6B";
								ro_addr_counter := ro_addr_counter + 1;
							when 105 =>
								s_addr_port_arr_i(2)<=x"6C";
								ro_addr_counter := ro_addr_counter + 1;
							when 106 =>
								s_addr_port_arr_i(2)<=x"6D";
								ro_addr_counter := ro_addr_counter + 1;
							when 107 =>
								s_addr_port_arr_i(2)<=x"6E";
								ro_addr_counter := ro_addr_counter + 1;
							when 108 =>
								s_addr_port_arr_i(2)<=x"6F";
								ro_addr_counter := ro_addr_counter + 1;
							when 109 =>
								s_addr_port_arr_i(2)<=x"70";
								ro_addr_counter := ro_addr_counter + 1;
							when 110 =>
								s_addr_port_arr_i(2)<=x"71";
								ro_addr_counter := ro_addr_counter + 1;
							when 111 =>
								s_addr_port_arr_i(2)<=x"72";
								ro_addr_counter := ro_addr_counter + 1;
							when 112 =>
								s_addr_port_arr_i(2)<=x"73";
								ro_addr_counter := ro_addr_counter + 1;
							when 113 =>
								s_addr_port_arr_i(2)<=x"74";
								ro_addr_counter := ro_addr_counter + 1;
							when 114 =>
								s_addr_port_arr_i(2)<=x"75";
								ro_addr_counter := ro_addr_counter + 1;
							when 115 =>
								s_addr_port_arr_i(2)<=x"76";
								ro_addr_counter := ro_addr_counter + 1;
							when 116 =>
								s_addr_port_arr_i(2)<=x"77";
								ro_addr_counter := ro_addr_counter + 1;
							when 117 =>
								s_addr_port_arr_i(2)<=x"78";
								ro_addr_counter := ro_addr_counter + 1;
							when 118 =>
								s_addr_port_arr_i(2)<=x"79";
								ro_addr_counter := ro_addr_counter + 1;
							when 119 =>
								s_addr_port_arr_i(2)<=x"7A";
								ro_addr_counter := ro_addr_counter + 1;
							when 120 =>
								s_addr_port_arr_i(2)<=x"7B";
								ro_addr_counter := ro_addr_counter + 1;
							when 121 =>
								s_addr_port_arr_i(2)<=x"7C";
								ro_addr_counter := ro_addr_counter + 1;
							when 122 =>
								s_addr_port_arr_i(2)<=x"7D";
								ro_addr_counter := ro_addr_counter + 1;
							when 123 =>
								s_addr_port_arr_i(2)<=x"7E";
								ro_addr_counter := ro_addr_counter + 1;
							when 124 =>
								s_addr_port_arr_i(2)<=x"7F";
								ro_addr_counter := ro_addr_counter + 1;
							when 125 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"8";  --Read enable on port a of ram 3
								s_addr_port_arr_i(3)<=x"00";
							when 126 =>
								ro_addr_counter := ro_addr_counter + 1;
								s3_pipe_rden_i<=x"8";  --Read enable on port a of ram 3
								s_addr_port_arr_i(3)<=x"01";
							when 127 =>
							ro_addr_counter := 0;
								s3_pipe_rden_i<=x"8";  --Read enable on port a of ram 3
								s_addr_port_arr_i(3)<=x"02";
								ram_counter:= ram_counter + 1; --Increment RAM counter
							when others =>
						end case;
					when 3 =>
						s3_pipe_rden_i<=x"8"; --Read enable on port a of ram 4
					   s3_pipeO.s3_pipe_data_o<=s_data_port_arr_o(3); --Direct output data to sub ram data out
						case ro_addr_counter is 
							when 0 =>
								s_addr_port_arr_i(3)<=x"03";
								ro_addr_counter := ro_addr_counter + 1;
							when 1 =>
								s_addr_port_arr_i(3)<=x"04";
								ro_addr_counter := ro_addr_counter + 1;
							when 2 =>
								s_addr_port_arr_i(3)<=x"05";
								ro_addr_counter := ro_addr_counter + 1;
							when 3 =>
								s_addr_port_arr_i(3)<=x"06";
								ro_addr_counter := ro_addr_counter + 1;
							when 4 =>
								s_addr_port_arr_i(3)<=x"07";
								ro_addr_counter := ro_addr_counter + 1;
							when 5 =>
								s_addr_port_arr_i(3)<=x"08";
								ro_addr_counter := ro_addr_counter + 1;
							when 6 =>
								s_addr_port_arr_i(3)<=x"09";
								ro_addr_counter := ro_addr_counter + 1;
							when 7 =>
								s_addr_port_arr_i(3)<=x"0A";
								ro_addr_counter := ro_addr_counter + 1;
							when 8 =>
								s_addr_port_arr_i(3)<=x"0B";
								ro_addr_counter := ro_addr_counter + 1;
							when 9 =>
								s_addr_port_arr_i(3)<=x"0C";
								ro_addr_counter := ro_addr_counter + 1;
							when 10 =>
								s_addr_port_arr_i(3)<=x"0D";
								ro_addr_counter := ro_addr_counter + 1;
							when 11 =>
								s_addr_port_arr_i(3)<=x"0E";
								ro_addr_counter := ro_addr_counter + 1;
							when 12 =>
								s_addr_port_arr_i(3)<=x"0F";
								ro_addr_counter := ro_addr_counter + 1;
							when 13 =>
								s_addr_port_arr_i(3)<=x"10";
								ro_addr_counter := ro_addr_counter + 1;
							when 14 =>
								s_addr_port_arr_i(3)<=x"11";
								ro_addr_counter := ro_addr_counter + 1;
							when 15 =>
								s_addr_port_arr_i(3)<=x"12";
								ro_addr_counter := ro_addr_counter + 1;
							when 16 =>
								s_addr_port_arr_i(3)<=x"13";
								ro_addr_counter := ro_addr_counter + 1;
							when 17 =>
								s_addr_port_arr_i(3)<=x"14";
								ro_addr_counter := ro_addr_counter + 1;
							when 18 =>
								s_addr_port_arr_i(3)<=x"15";
								ro_addr_counter := ro_addr_counter + 1;
							when 19 =>
								s_addr_port_arr_i(3)<=x"16";
								ro_addr_counter := ro_addr_counter + 1;
							when 20 =>
								s_addr_port_arr_i(3)<=x"17";
								ro_addr_counter := ro_addr_counter + 1;
							when 21 =>
								s_addr_port_arr_i(3)<=x"18";
								ro_addr_counter := ro_addr_counter + 1;
							when 22 =>
								s_addr_port_arr_i(3)<=x"19";
								ro_addr_counter := ro_addr_counter + 1;
							when 23 =>
								s_addr_port_arr_i(3)<=x"1A";
								ro_addr_counter := ro_addr_counter + 1;
							when 24 =>
								s_addr_port_arr_i(3)<=x"1B";
								ro_addr_counter := ro_addr_counter + 1;
							when 25 =>
								s_addr_port_arr_i(3)<=x"1C";
								ro_addr_counter := ro_addr_counter + 1;
							when 26 =>
								s_addr_port_arr_i(3)<=x"1D";
								ro_addr_counter := ro_addr_counter + 1;
							when 27 =>
								s_addr_port_arr_i(3)<=x"1E";
								ro_addr_counter := ro_addr_counter + 1;
							when 28 =>
								s_addr_port_arr_i(3)<=x"1F";
								ro_addr_counter := ro_addr_counter + 1;
							when 29 =>
								s_addr_port_arr_i(3)<=x"20";
								ro_addr_counter := ro_addr_counter + 1;
							when 30 =>
								s_addr_port_arr_i(3)<=x"21";
								ro_addr_counter := ro_addr_counter + 1;
							when 31 =>
								s_addr_port_arr_i(3)<=x"22";
								ro_addr_counter := ro_addr_counter + 1;
							when 32 =>
								s_addr_port_arr_i(3)<=x"23";
								ro_addr_counter := ro_addr_counter + 1;
							when 33 =>
								s_addr_port_arr_i(3)<=x"24";
								ro_addr_counter := ro_addr_counter + 1;
							when 34 =>
								s_addr_port_arr_i(3)<=x"25";
								ro_addr_counter := ro_addr_counter + 1;
							when 35 =>
								s_addr_port_arr_i(3)<=x"26";
								ro_addr_counter := ro_addr_counter + 1;
							when 36 =>
								s_addr_port_arr_i(3)<=x"27";
								ro_addr_counter := ro_addr_counter + 1;
							when 37 =>
								s_addr_port_arr_i(3)<=x"28";
								ro_addr_counter := ro_addr_counter + 1;
							when 38 =>
								s_addr_port_arr_i(3)<=x"29";
								ro_addr_counter := ro_addr_counter + 1;
							when 39 =>
								s_addr_port_arr_i(3)<=x"2A";
								ro_addr_counter := ro_addr_counter + 1;
							when 40 =>
								s_addr_port_arr_i(3)<=x"2B";
								ro_addr_counter := ro_addr_counter + 1;
							when 41 =>
								s_addr_port_arr_i(3)<=x"2C";
								ro_addr_counter := ro_addr_counter + 1;
							when 42 =>
								s_addr_port_arr_i(3)<=x"2D";
								ro_addr_counter := ro_addr_counter + 1;
							when 43 =>
								s_addr_port_arr_i(3)<=x"2E";
								ro_addr_counter := ro_addr_counter + 1;
							when 44 =>
								s_addr_port_arr_i(3)<=x"2F";
								ro_addr_counter := ro_addr_counter + 1;
							when 45 =>
								s_addr_port_arr_i(3)<=x"30";
								ro_addr_counter := ro_addr_counter + 1;
							when 46 =>
								s_addr_port_arr_i(3)<=x"31";
								ro_addr_counter := ro_addr_counter + 1;
							when 47 =>
								s_addr_port_arr_i(3)<=x"32";
								ro_addr_counter := ro_addr_counter + 1;
							when 48 =>
								s_addr_port_arr_i(3)<=x"33";
								ro_addr_counter := ro_addr_counter + 1;
							when 49 =>
								s_addr_port_arr_i(3)<=x"34";
								ro_addr_counter := ro_addr_counter + 1;
							when 50 =>
								s_addr_port_arr_i(3)<=x"35";
								ro_addr_counter := ro_addr_counter + 1;
							when 51 =>
								s_addr_port_arr_i(3)<=x"36";
								ro_addr_counter := ro_addr_counter + 1;
							when 52 =>
								s_addr_port_arr_i(3)<=x"37";
								ro_addr_counter := ro_addr_counter + 1;
							when 53 =>
								s_addr_port_arr_i(3)<=x"38";
								ro_addr_counter := ro_addr_counter + 1;
							when 54 =>
								s_addr_port_arr_i(3)<=x"39";
								ro_addr_counter := ro_addr_counter + 1;
							when 55 =>
								s_addr_port_arr_i(3)<=x"3A";
								ro_addr_counter := ro_addr_counter + 1;
							when 56 =>
								s_addr_port_arr_i(3)<=x"3B";
								ro_addr_counter := ro_addr_counter + 1;
							when 57 =>
								s_addr_port_arr_i(3)<=x"3C";
								ro_addr_counter := ro_addr_counter + 1;
							when 58 =>
								s_addr_port_arr_i(3)<=x"3D";
								ro_addr_counter := ro_addr_counter + 1;
							when 59 =>
								s_addr_port_arr_i(3)<=x"3E";
								ro_addr_counter := ro_addr_counter + 1;
							when 60 =>
								s_addr_port_arr_i(3)<=x"3F";
								ro_addr_counter := ro_addr_counter + 1;
							when 61 =>
								s_addr_port_arr_i(3)<=x"40";
								ro_addr_counter := ro_addr_counter + 1;
							when 62 =>
								s_addr_port_arr_i(3)<=x"41";
								ro_addr_counter := ro_addr_counter + 1;
							when 63 =>
								s_addr_port_arr_i(3)<=x"42";
								ro_addr_counter := ro_addr_counter + 1;
							when 64 =>
								s_addr_port_arr_i(3)<=x"43";
								ro_addr_counter := ro_addr_counter + 1;
							when 65 =>
								s_addr_port_arr_i(3)<=x"44";
								ro_addr_counter := ro_addr_counter + 1;
							when 66 =>
								s_addr_port_arr_i(3)<=x"45";
								ro_addr_counter := ro_addr_counter + 1;
							when 67 =>
								s_addr_port_arr_i(3)<=x"46";
								ro_addr_counter := ro_addr_counter + 1;
							when 68 =>
								s_addr_port_arr_i(3)<=x"47";
								ro_addr_counter := ro_addr_counter + 1;
							when 69 =>
								s_addr_port_arr_i(3)<=x"48";
								ro_addr_counter := ro_addr_counter + 1;
							when 70 =>
								s_addr_port_arr_i(3)<=x"49";
								ro_addr_counter := ro_addr_counter + 1;
							when 71 =>
								s_addr_port_arr_i(3)<=x"4A";
								ro_addr_counter := ro_addr_counter + 1;
							when 72 =>
								s_addr_port_arr_i(3)<=x"4B";
								ro_addr_counter := ro_addr_counter + 1;
							when 73 =>
								s_addr_port_arr_i(3)<=x"4C";
								ro_addr_counter := ro_addr_counter + 1;
							when 74 =>
								s_addr_port_arr_i(3)<=x"4D";
								ro_addr_counter := ro_addr_counter + 1;
							when 75 =>
								s_addr_port_arr_i(3)<=x"4E";
								ro_addr_counter := ro_addr_counter + 1;
							when 76 =>
								s_addr_port_arr_i(3)<=x"4F";
								ro_addr_counter := ro_addr_counter + 1;
							when 77 =>
								s_addr_port_arr_i(3)<=x"50";
								ro_addr_counter := ro_addr_counter + 1;
							when 78 =>
								s_addr_port_arr_i(3)<=x"51";
								ro_addr_counter := ro_addr_counter + 1;
							when 79 =>
								s_addr_port_arr_i(3)<=x"52";
								ro_addr_counter := ro_addr_counter + 1;
							when 80 =>
								s_addr_port_arr_i(3)<=x"53";
								ro_addr_counter := ro_addr_counter + 1;
							when 81 =>
								s_addr_port_arr_i(3)<=x"54";
								ro_addr_counter := ro_addr_counter + 1;
							when 82 =>
								s_addr_port_arr_i(3)<=x"55";
								ro_addr_counter := ro_addr_counter + 1;
							when 83 =>
								s_addr_port_arr_i(3)<=x"56";
								ro_addr_counter := ro_addr_counter + 1;
							when 84 =>
								s_addr_port_arr_i(3)<=x"57";
								ro_addr_counter := ro_addr_counter + 1;
							when 85 =>
								s_addr_port_arr_i(3)<=x"58";
								ro_addr_counter := ro_addr_counter + 1;
							when 86 =>
								s_addr_port_arr_i(3)<=x"59";
								ro_addr_counter := ro_addr_counter + 1;
							when 87 =>
								s_addr_port_arr_i(3)<=x"5A";
								ro_addr_counter := ro_addr_counter + 1;
							when 88 =>
								s_addr_port_arr_i(3)<=x"5B";
								ro_addr_counter := ro_addr_counter + 1;
							when 89 =>
								s_addr_port_arr_i(3)<=x"5C";
								ro_addr_counter := ro_addr_counter + 1;
							when 90 =>
								s_addr_port_arr_i(3)<=x"5D";
								ro_addr_counter := ro_addr_counter + 1;
							when 91 =>
								s_addr_port_arr_i(3)<=x"5E";
								ro_addr_counter := ro_addr_counter + 1;
							when 92 =>
								s_addr_port_arr_i(3)<=x"5F";
								ro_addr_counter := ro_addr_counter + 1;
							when 93 =>
								s_addr_port_arr_i(3)<=x"60";
								ro_addr_counter := ro_addr_counter + 1;
							when 94 =>
								s_addr_port_arr_i(3)<=x"61";
								ro_addr_counter := ro_addr_counter + 1;
							when 95 =>
								s_addr_port_arr_i(3)<=x"62";
								ro_addr_counter := ro_addr_counter + 1;
							when 96 =>
								s_addr_port_arr_i(3)<=x"63";
								ro_addr_counter := ro_addr_counter + 1;
							when 97 =>
								s_addr_port_arr_i(3)<=x"64";
								ro_addr_counter := ro_addr_counter + 1;
							when 98 =>
								s_addr_port_arr_i(3)<=x"65";
								ro_addr_counter := ro_addr_counter + 1;
							when 99 =>
								s_addr_port_arr_i(3)<=x"66";
								ro_addr_counter := ro_addr_counter + 1;
							when 100 =>
								s_addr_port_arr_i(3)<=x"67";
								ro_addr_counter := ro_addr_counter + 1;
							when 101 =>
								s_addr_port_arr_i(3)<=x"68";
								ro_addr_counter := ro_addr_counter + 1;
							when 102 =>
								s_addr_port_arr_i(3)<=x"69";
								ro_addr_counter := ro_addr_counter + 1;
							when 103 =>
								s_addr_port_arr_i(3)<=x"6A";
								ro_addr_counter := ro_addr_counter + 1;
							when 104 =>
								s_addr_port_arr_i(3)<=x"6B";
								ro_addr_counter := ro_addr_counter + 1;
							when 105 =>
								s_addr_port_arr_i(3)<=x"6C";
								ro_addr_counter := ro_addr_counter + 1;
							when 106 =>
								s_addr_port_arr_i(3)<=x"6D";
								ro_addr_counter := ro_addr_counter + 1;
							when 107 =>
								s_addr_port_arr_i(3)<=x"6E";
								ro_addr_counter := ro_addr_counter + 1;
							when 108 =>
								s_addr_port_arr_i(3)<=x"6F";
								ro_addr_counter := ro_addr_counter + 1;
							when 109 =>
								s_addr_port_arr_i(3)<=x"70";
								ro_addr_counter := ro_addr_counter + 1;
							when 110 =>
								s_addr_port_arr_i(3)<=x"71";
								ro_addr_counter := ro_addr_counter + 1;
							when 111 =>
								s_addr_port_arr_i(3)<=x"72";
								ro_addr_counter := ro_addr_counter + 1;
							when 112 =>
								s_addr_port_arr_i(3)<=x"73";
								ro_addr_counter := ro_addr_counter + 1;
							when 113 =>
								s_addr_port_arr_i(3)<=x"74";
								ro_addr_counter := ro_addr_counter + 1;
							when 114 =>
								s_addr_port_arr_i(3)<=x"75";
								ro_addr_counter := ro_addr_counter + 1;
							when 115 =>
								s_addr_port_arr_i(3)<=x"76";
								ro_addr_counter := ro_addr_counter + 1;
							when 116 =>
								s_addr_port_arr_i(3)<=x"77";
								ro_addr_counter := ro_addr_counter + 1;
							when 117 =>
								s_addr_port_arr_i(3)<=x"78";
								ro_addr_counter := ro_addr_counter + 1;
							when 118 =>
								s_addr_port_arr_i(3)<=x"79";
								ro_addr_counter := ro_addr_counter + 1;
							when 119 =>
								s_addr_port_arr_i(3)<=x"7A";
								ro_addr_counter := ro_addr_counter + 1;
							when 120 =>
								s_addr_port_arr_i(3)<=x"7B";
								ro_addr_counter := ro_addr_counter + 1;
							when 121 =>
								s_addr_port_arr_i(3)<=x"7C";
								ro_addr_counter := ro_addr_counter + 1;
							when 122 =>
								s_addr_port_arr_i(3)<=x"7D";
								ro_addr_counter := ro_addr_counter + 1;
							when 123 =>
								s_addr_port_arr_i(3)<=x"7E";
								ro_addr_counter := ro_addr_counter + 1;
							when 124 =>
								s_addr_port_arr_i(3)<=x"7F";
								ro_addr_counter := ro_addr_counter + 1;
							when 125 =>
								ro_addr_counter := ro_addr_counter + 1;
							when 126 =>
								ro_addr_counter := ro_addr_counter + 1;
							when 127 =>
								ro_addr_counter := ro_addr_counter + 1;
							when 128 =>
								s3_pipeO.s3_pipe_data_v_o<='0';
								s3_pipe_rden_i<=x"0";
								ro_addr_counter := 0;
							when others =>
						end case;
					when others =>
				end case;
			end if;
		end if;
	end process;	
			
end main;